module circuit(x, y);
  // x is the input
  // y is the output
  // Good luck and have fun
  wire admiringbardeen;
  wire admiringhelga;
  wire admiringride;
  wire adoringbassi;
  wire adoringbohr;
  wire adoringdhawan;
  wire adoringhook;
  wire adoringmargulis;
  wire affectionatebell;
  wire affectionatehazel;
  wire agitatedbose;
  wire agitatedharold;
  wire amazinghiro;
  wire amazingkermit;
  wire amazingmclean;
  wire amazingshaw;
  wire angrywozniak;
  wire awesomegauss;
  wire awesomeheisenberg;
  wire beautifuldarwin;
  wire blissfulalbattani;
  wire blissfulheihei;
  wire blissfulnewton;
  wire boldishizaka;
  wire boringheyrovsky;
  wire bravehoney;
  wire braveivan;
  wire bravekata;
  wire busyjoliot;
  wire busynorthcutt;
  wire charmingjunior;
  wire compassionatecray;
  wire compassionatehiram;
  wire compassionatejose;
  wire competentaustin;
  wire competenthatbox;
  wire competentichabod;
  wire competentwilliamson;
  wire condescendingsatoshi;
  wire confidentagnesi;
  wire confidentbouman;
  wire cooljackjack;
  wire coolkc;
  wire crankykeldysh;
  wire crazycarson;
  wire dazzlingcannon;
  wire dazzlingjerry;
  wire dazzlingjudge;
  wire determinedcartwright;
  wire determinedgus;
  wire determinedinaki;
  wire dreamygustavo;
  wire eagerkare;
  wire eagerkilby;
  wire eagerpoincare;
  wire ecstaticbuck;
  wire ecstaticshockley;
  wire ecstaticsinoussi;
  wire elasticborg;
  wire elasticburnell;
  wire elasticiago;
  wire elasticjill;
  wire elatedharper;
  wire elatedhedgie;
  wire elegantblack;
  wire elegantdavinci;
  wire elegantkaa;
  wire elegantmerkle;
  wire eloquentkaren;
  wire excitingcarver;
  wire excitingcerf;
  wire excitinghoonah;
  wire excitingjackson;
  wire excitingjesse;
  wire ferventjeb;
  wire ferventjin;
  wire festivechandrasekhar;
  wire festivegrothendieck;
  wire festiveperlman;
  wire flamboyantchatelet;
  wire flamboyantleavitt;
  wire focusedgalileo;
  wire focusedjepsen;
  wire focusedshamir;
  wire friendlyhamilton;
  wire friendlyharry;
  wire friendlyjenny;
  wire frostyjasmine;
  wire frostyjennings;
  wire frostyswanson;
  wire frostyvolhard;
  wire funnygoldwasser;
  wire funnyleakey;
  wire funnyshtern;
  wire gallanthellman;
  wire gallantmirzakhani;
  wire giftedgoodall;
  wire giftedwilson;
  wire goofychebyshev;
  wire goofyjunia;
  wire goofysammet;
  wire goofystonebraker;
  wire graciousgermain;
  wire graciousherb;
  wire graciousknuth;
  wire greatelbakyan;
  wire greatjames;
  wire greatmoser;
  wire happybrahmagupta;
  wire happydriscoll;
  wire hardcorecurie;
  wire hardcorejuanita;
  wire hardcorejulio;
  wire hardcorerubin;
  wire heuristicchaum;
  wire heuristicgagarin;
  wire heuristichaslett;
  wire hopefulhaibt;
  wire hopefulkele;
  wire hungryjane;
  wire hungrynash;
  wire hungrywright;
  wire hungryzhukovsky;
  wire infallibleblackwell;
  wire infalliblegolick;
  wire infalliblejake;
  wire infalliblejason;
  wire infalliblejoy;
  wire inspiringfermi;
  wire inspiringisabela;
  wire inspiringjang;
  wire inspiringjiminy;
  wire intelligenthermes;
  wire intelligentnoether;
  wire interestingeuclid;
  wire interestinghawking;
  wire interestinglamport;
  wire jollyedison;
  wire jollyjorge;
  wire jovialgoldberg;
  wire jovialgyro;
  wire jovialhenrietta;
  wire jovialhera;
  wire jovialhoneymaren;
  wire joviallehmann;
  wire jovialwiles;
  wire kindhector;
  wire kindherschel;
  wire kindrosalind;
  wire laughingalmeida;
  wire laughingbhaskara;
  wire laughingdubinsky;
  wire laughingmccarthy;
  wire laughingmorse;
  wire laughingsaha;
  wire lovingdirac;
  wire lovingeasley;
  wire lovinghoagy;
  wire lovingjemison;
  wire lovingkowalevski;
  wire lovingmoore;
  wire lucidbabbage;
  wire lucidjaeger;
  wire lucidpike;
  wire lucidsolomon;
  wire magicalchaplygin;
  wire magicaljudy;
  wire magicalken;
  wire magicalliskov;
  wire magicalwescoff;
  wire modestfeynman;
  wire modestjelly;
  wire modestmontalcini;
  wire modestshirley;
  wire modestswartz;
  wire modestvillani;
  wire musingholley;
  wire mystifyingbartik;
  wire mystifyinggates;
  wire naughtybooth;
  wire naughtyjangles;
  wire naughtynapier;
  wire nervoushonker;
  wire nervousmatsumoto;
  wire nervoustharp;
  wire nervousvisvesvaraya;
  wire niceclarke;
  wire nicefermat;
  wire niceganguly;
  wire nicejoshamee;
  wire niftyian;
  wire niftysnyder;
  wire nostalgicbrattain;
  wire nostalgiccori;
  wire nostalgichannah;
  wire objectivedijkstra;
  wire objectivejones;
  wire objectivelewin;
  wire objectivespence;
  wire optimisticptolemy;
  wire optimisticvarahamihira;
  wire peacefulardinghelli;
  wire peacefulsutherland;
  wire peacefulhermann;
  wire peacefuljackson;
  wire peacefulwing;
  wire pedanticcurran;
  wire pedantichumbert;
  wire pedantickari;
  wire pedantickhayyam;
  wire pedanticmeninsky;
  wire pedanticmurdock;
  wire pensivehailey;
  wire pensivemendeleev;
  wire practicaljubileena;
  wire practicalpayne;
  wire pricelesskalam;
  wire pricelesskevin;
  wire pricelessmeitner;
  wire quirkylederberg;
  wire quirkymendel;
  wire quirkyyalow;
  wire quizzicalhertz;
  wire quizzicalhugo;
  wire quizzicaljacques;
  wire quizzicalkala;
  wire quizzicalneumann;
  wire quizzicalpanini;
  wire recursinghallie;
  wire recursingraman;
  wire relaxedvaughan;
  wire reverentjohn;
  wire reverentjonah;
  wire reverentroentgen;
  wire romantickapitsa;
  wire sadgould;
  wire sadjimmy;
  wire serenehissy;
  wire serenehofstadter;
  wire serenemahavira;
  wire sereneyonath;
  wire sharpheffalump;
  wire sharpnightingale;
  wire sharpproskuriakova;
  wire sillykekata;
  wire sleepygypsy;
  wire stoicelion;
  wire stoicfaraday;
  wire stoicgalois;
  wire stoichercules;
  wire stoickepler;
  wire stoicmcclintock;
  wire strangeelgamal;
  wire strangehappy;
  wire strangekhorana;
  wire stupefiedblackburn;
  wire stupefiedhopper;
  wire stupefiedjiku;
  wire stupefiedjohnnie;
  wire suspiciousjim;
  wire sweetcryptanalyse;
  wire sweetimelda;
  wire sweetinnoko;
  wire tenderallen;
  wire tenderellis;
  wire tenderfranklin;
  wire tendermestorf;
  wire thirstychatterjee;
  wire thirstygusto;
  wire thirstymclaren;
  wire trustingcolden;
  wire trustinghades;
  wire trustingtesla;
  wire unruffledgwen;
  wire unruffledhenry;
  wire unruffledhoover;
  wire unruffledhudson;
  wire unruffledkatie;
  wire unruffledsanderson;
  wire unruffledswirles;
  wire upbeatbanzai;
  wire upbeathurley;
  wire vibranthodgkin;
  wire vibranthorace;
  wire vigoroushit;
  wire wizardlylichterman;
  wire wonderfulboyd;
  wire wonderfulrobinson;
  wire xenodochialjack;
  wire xenodochiallumiere;
  wire xenodochialwilliams;
  wire youthfulantonelli;
  wire youthfularyabhata;
  wire youthfulturing;
  wire zealouslovelace;
  wire zealoustorvalds;
  wire zenbanach;
  wire zenhypatia;
  wire zenritchie;
  input [15:0] x;
  wire [15:0] x;
  output [15:0] y;
  wire [15:0] y;
  NAND admiringbell (.A(lovingkowalevski), .B(angrywozniak), .Y(happydriscoll));
  NAND adoringjames (.A(stoickepler), .B(reverentjohn), .Y(dazzlingjerry));
  NAND adoringstonebraker (.A(jovialgoldberg), .B(elasticiago), .Y(hungrywright));
  NAND blissfultaussig (.A(sweetimelda), .B(eagerpoincare), .Y(trustingcolden));
  NAND cleverkare (.A(competentichabod), .B(quirkymendel), .Y(goofysammet));
  NAND cleverpayne (.A(hungrynash), .B(pedanticmeninsky), .Y(greatelbakyan));
  NAND dazzlingkanga (.A(flamboyantleavitt), .B(kindherschel), .Y(awesomeheisenberg));
  NAND elegantrhodes (.A(pedantickhayyam), .B(heuristicchaum), .Y(upbeatbanzai));
  NAND festiveswartz (.A(elatedharper), .B(sadgould), .Y(joviallehmann));
  NAND flamboyantjill (.A(funnygoldwasser), .B(frostyvolhard), .Y(naughtyjangles));
  NAND greatbooth (.A(modestshirley), .B(focusedshamir), .Y(nervousmatsumoto));
  NAND happyheimlich (.A(compassionatejose), .B(magicalken), .Y(stoicfaraday));
  NAND intelligentcartwright (.A(jollyjorge), .B(niceganguly), .Y(elegantdavinci));
  NAND interestingjessie (.A(youthfulantonelli), .B(blissfulalbattani), .Y(braveivan));
  NAND lovingeinstein (.A(quizzicalpanini), .B(hardcorecurie), .Y(magicalliskov));
  NAND niftyrobinson (.A(infalliblejason), .B(zealoustorvalds), .Y(goofyjunia));
  NAND optimisticjustin (.A(kindhector), .B(peacefulhermann), .Y(peacefuljackson));
  NAND sadhypatia (.A(agitatedharold), .B(thirstygusto), .Y(excitingcerf));
  NAND suspiciousdewdney (.A(heuristicgagarin), .B(lovingmoore), .Y(tenderfranklin));
  NAND xenodochialbenz (.A(crankykeldysh), .B(sleepygypsy), .Y(youthfularyabhata));
  NOR cleverkelsi (.A(quizzicalpanini), .B(tenderallen), .Y(hardcorejulio));
  NOR ecstaticwescoff (.A(frostyvolhard), .B(coolkc), .Y(eloquentkaren));
  NOR eloquentvaughan (.A(zealoustorvalds), .B(tenderellis), .Y(laughingbhaskara));
  NOR excitingjennings (.A(xenodochiallumiere), .B(trustingtesla), .Y(goofychebyshev));
  NOR ferventhamm (.A(blissfulalbattani), .B(heuristicchaum), .Y(inspiringjiminy));
  NOR flamboyantbeaver (.A(hardcorecurie), .B(heuristicgagarin), .Y(adoringhook));
  NOR frostyharv (.A(festiveperlman), .B(infalliblejason), .Y(admiringbardeen));
  NOR frostyhit (.A(peacefulhermann), .B(stoicmcclintock), .Y(hardcorejuanita));
  NOR hardcorejennifer (.A(magicalken), .B(jollyjorge), .Y(infalliblegolick));
  NOR hardcorenobel (.A(lovingjemison), .B(adoringbohr), .Y(elegantmerkle));
  NOR heuristicfeynman (.A(peacefulardinghelli), .B(wizardlylichterman), .Y(lucidpike));
  NOR heuristichank (.A(youthfulantonelli), .B(sweetimelda), .Y(sadjimmy));
  NOR intelligenttu (.A(kindherschel), .B(stoicgalois), .Y(amazingkermit));
  NOR interestingchaplygin (.A(quirkymendel), .B(hungrynash), .Y(hungryzhukovsky));
  NOR interestingjack (.A(elasticiago), .B(agitatedharold), .Y(funnyleakey));
  NOR magicalsutherland (.A(pricelesskevin), .B(pedanticmeninsky), .Y(cooljackjack));
  NOR magicalhonker (.A(friendlyjenny), .B(jovialgoldberg), .Y(mystifyinggates));
  NOR modesthopper (.A(nostalgicbrattain), .B(elatedharper), .Y(mystifyingbartik));
  NOR modestnoyce (.A(interestinglamport), .B(confidentbouman), .Y(pedantickari));
  NOR modestsolomon (.A(kindrosalind), .B(modestvillani), .Y(sereneyonath));
  NOR nostalgicjuarez (.A(eagerpoincare), .B(crankykeldysh), .Y(interestinghawking));
  NOR objectivefermi (.A(dazzlingjudge), .B(focusedshamir), .Y(stupefiedjohnnie));
  NOR relaxedhamster (.A(kindhector), .B(stoickepler), .Y(adoringbassi));
  NOR thirstyroentgen (.A(competentichabod), .B(sadgould), .Y(amazingshaw));
  NOR trustingarchimedes (.A(compassionatehiram), .B(angrywozniak), .Y(practicaljubileena));
  NOR wizardlycurran (.A(unruffledswirles), .B(thirstygusto), .Y(affectionatehazel));
  NOR youthfulhuey (.A(sleepygypsy), .B(unruffledhudson), .Y(elegantblack));
  NOT agitatedizzy (.A(sleepygypsy), .Y(pedantickhayyam));
  NOT condescendingjoe (.A(blissfulalbattani), .Y(trustinghades));
  NOT greatlalande (.A(sweetimelda), .Y(interestinglamport));
  NOT quirkyptolemy (.A(competentichabod), .Y(elegantkaa));
  NOT youtu_be (.A(heuristicchaum), .Y(unruffledhudson));
  NOT pJMH1Oye8f8 (.A(hungrynash), .Y(dreamygustavo));
  NOT trustingian (.A(nostalgicbrattain), .Y(pricelesskevin));
  NOT trustingramanujan (.A(eagerpoincare), .Y(confidentbouman));
  XOR adoringbuck (.A(reverentjohn), .B(sharpnightingale), .Y(thirstygusto));
  XOR adoringhissy (.A(dazzlingjerry), .B(nervoustharp), .Y(elasticiago));
  XOR adoringjonah (.A(elegantdavinci), .B(excitingcarver), .Y(funnygoldwasser));
  XOR angrycohen (.A(naughtynapier), .B(inspiringjiminy), .Y(vibranthodgkin));
  XOR awesomehera (.A(nervousmatsumoto), .B(bravekata), .Y(stoicelion));
  XOR awesomekate (.A(pedantickari), .B(pensivehailey), .Y(zealoustorvalds));
  XOR beautifulheyrovsky (.A(niceganguly), .B(quirkyyalow), .Y(modestvillani));
  XOR blissfulhaslett (.A(funnyleakey), .B(bravehoney), .Y(elatedharper));
  XOR blissfulhoneymaren (.A(tenderallen), .B(stupefiedjohnnie), .Y(quirkyyalow));
  XOR blissfulnorthcutt (.A(compassionatehiram), .B(stupefiedjohnnie), .Y(flamboyantchatelet));
  XOR boldeuler (.A(youthfulantonelli), .B(agitatedbose), .Y(pensivehailey));
  XOR boringgoldstine (.A(elegantmerkle), .B(elatedhedgie), .Y(compassionatejose));
  XOR boringlamarr (.A(lucidjaeger), .B(hardcorejulio), .Y(magicalken));
  XOR boringmargulis (.A(peacefulhermann), .B(funnyleakey), .Y(zenritchie));
  XOR bravejock (.A(tenderfranklin), .B(ferventjeb), .Y(stoicgalois));
  XOR busykenai (.A(sadjimmy), .B(festivegrothendieck), .Y(angrywozniak));
  XOR cleverjohnny (.A(agitatedbose), .B(trustingcolden), .Y(ferventjeb));
  XOR cleverjohnson (.A(confidentbouman), .B(elegantmerkle), .Y(dazzlingcannon));
  XOR compassionatesaha (.A(sharpnightingale), .B(goofychebyshev), .Y(quirkymendel));
  XOR competentbanach (.A(funnygoldwasser), .B(sharpnightingale), .Y(objectivedijkstra));
  XOR competenthelga (.A(tendermestorf), .B(lucidpike), .Y(hungrynash));
  XOR condescendingpare (.A(admiringbardeen), .B(ferventjeb), .Y(dazzlingjudge));
  XOR confidenthopper (.A(sadjimmy), .B(inspiringisabela), .Y(tenderellis));
  XOR confidentkapitsa (.A(adoringbassi), .B(magicaljudy), .Y(jovialgoldberg));
  XOR dazzlingmendeleev (.A(crankykeldysh), .B(hardcorejulio), .Y(competentaustin));
  XOR eagerlewin (.A(flamboyantchatelet), .B(hardcorejuanita), .Y(wizardlylichterman));
  XOR elatedbhabha (.A(peacefuljackson), .B(friendlyhamilton), .Y(peacefulardinghelli));
  XOR elatedjessica (.A(sweetimelda), .B(strangekhorana), .Y(infalliblejason));
  XOR elegantburnell (.A(stoicelion), .B(tendermestorf), .Y(unruffledswirles));
  XOR epicdhawan (.A(nervousmatsumoto), .B(modestmontalcini), .Y(frostyvolhard));
  XOR epicjane (.A(modestjelly), .B(happydriscoll), .Y(modestshirley));
  XOR festivewu (.A(interestinglamport), .B(adoringhook), .Y(intelligentnoether));
  XOR friendlygreider (.A(angrywozniak), .B(amazingkermit), .Y(frostyjasmine));
  XOR frostyhitchhiking (.A(awesomeheisenberg), .B(laughingmccarthy), .Y(peacefulhermann));
  XOR funnyjafar (.A(crankykeldysh), .B(youthfulturing), .Y(recursingraman));
  XOR gallanthatbox (.A(excitingcerf), .B(condescendingsatoshi), .Y(sadgould));
  XOR hardcorehugle (.A(elegantblack), .B(recursingraman), .Y(adoringbohr));
  XOR heuristichertz (.A(amazingkermit), .B(nostalgiccori), .Y(stoicmcclintock));
  XOR heuristickeller (.A(pedantickhayyam), .B(vibranthodgkin), .Y(lovingjemison));
  XOR hopefuljuan (.A(awesomeheisenberg), .B(lovingkowalevski), .Y(magicaljudy));
  XOR intelligentagnesi (.A(jollyjorge), .B(sereneyonath), .Y(tendermestorf));
  XOR intelligentblackburn (.A(blissfulalbattani), .B(goofyjunia), .Y(nostalgiccori));
  XOR intelligentmclaren (.A(frostyvolhard), .B(tendermestorf), .Y(xenodochiallumiere));
  XOR interestinghenry (.A(naughtyjangles), .B(sweetinnoko), .Y(agitatedharold));
  XOR interestingmurdock (.A(trustinghades), .B(goofyjunia), .Y(serenemahavira));
  XOR jollycray (.A(modestshirley), .B(hardcorejuanita), .Y(stupefiedjiku));
  XOR jollyneumann (.A(friendlyjenny), .B(boldishizaka), .Y(nostalgicbrattain));
  XOR jollyproskuriakova (.A(magicalken), .B(eloquentkaren), .Y(sharpnightingale));
  XOR keenmayer (.A(unruffledhudson), .B(modestjelly), .Y(tenderallen));
  XOR kindkele (.A(quirkyyalow), .B(hardcorejuanita), .Y(trustingtesla));
  XOR kindwing (.A(hungrywright), .B(kindrosalind), .Y(boldishizaka));
  XOR laughingjepsen (.A(heuristicgagarin), .B(infalliblegolick), .Y(sweetinnoko));
  XOR laughingwiles (.A(modestjelly), .B(laughingbhaskara), .Y(niceganguly));
  XOR lucidjeff (.A(youthfularyabhata), .B(excitingjackson), .Y(heuristicgagarin));
  XOR magicalgauss (.A(hardcorecurie), .B(magicalken), .Y(excitingcarver));
  XOR magicalhorace (.A(modestshirley), .B(quirkyyalow), .Y(coolkc));
  XOR modestharley (.A(unruffledgwen), .B(braveivan), .Y(modestjelly));
  XOR modestkirch (.A(infalliblejoy), .B(interestinghawking), .Y(strangekhorana));
  XOR musingdiffie (.A(interestinglamport), .B(strangekhorana), .Y(lovingmoore));
  XOR mystifyingjake (.A(amazingkermit), .B(serenemahavira), .Y(kindrosalind));
  XOR mystifyingmaxwell (.A(youthfularyabhata), .B(pricelesskalam), .Y(festiveperlman));
  XOR naughtypascal (.A(blissfulalbattani), .B(optimisticvarahamihira), .Y(festivegrothendieck));
  XOR nervousbrown (.A(youthfulturing), .B(elegantblack), .Y(lucidjaeger));
  XOR nervousjett (.A(vibranthodgkin), .B(practicaljubileena), .Y(jollyjorge));
  XOR nicebabbage (.A(stoickepler), .B(affectionatehazel), .Y(lovingeasley));
  XOR nicejackal (.A(upbeatbanzai), .B(recursingraman), .Y(hardcorecurie));
  XOR nostalgicpasteur (.A(infalliblegolick), .B(dazzlingcannon), .Y(stoickepler));
  XOR optimisticcarson (.A(coolkc), .B(mystifyinggates), .Y(serenehofstadter));
  XOR optimistichappy (.A(goofyjunia), .B(jovialhenrietta), .Y(focusedshamir));
  XOR optimisticjang (.A(stoicfaraday), .B(infalliblejason), .Y(nervoustharp));
  XOR pedanticheadless (.A(magicalliskov), .B(elatedhedgie), .Y(flamboyantleavitt));
  XOR pensiveboyd (.A(objectivedijkstra), .B(greatelbakyan), .Y(funnyshtern));
  XOR practicalhoagy (.A(sleepygypsy), .B(practicaljubileena), .Y(bravekata));
  XOR pricelesskala (.A(stoicelion), .B(lucidpike), .Y(pedantichumbert));
  XOR pricelessthompson (.A(heuristicchaum), .B(modestjelly), .Y(compassionatehiram));
  XOR quizzicalchandrasekhar (.A(amazingshaw), .B(zenritchie), .Y(elasticborg));
  XOR relaxedgus (.A(dazzlingjudge), .B(adoringbassi), .Y(bravehoney));
  XOR relaxedhiro (.A(quirkymendel), .B(funnyshtern), .Y(jovialgyro));
  XOR romanticengelbart (.A(eagerpoincare), .B(ecstaticsinoussi), .Y(excitingjackson));
  XOR romanticmirzakhani (.A(kindhector), .B(excitingcerf), .Y(blissfulheihei));
  XOR sadmeitner (.A(mystifyinggates), .B(stupefiedjiku), .Y(pedanticmeninsky));
  XOR sadspence (.A(goofysammet), .B(blissfulheihei), .Y(hopefulhaibt));
  XOR serenemcnulty (.A(youthfulantonelli), .B(admiringbardeen), .Y(laughingmccarthy));
  XOR sillychatterjee (.A(affectionatehazel), .B(greatmoser), .Y(competentichabod));
  XOR sillyhannah (.A(mystifyingbartik), .B(serenehofstadter), .Y(sharpheffalump));
  XOR sillyjune (.A(stoicfaraday), .B(intelligentnoether), .Y(kindhector));
  XOR strangehellman (.A(hungryzhukovsky), .B(lovingeasley), .Y(nicejoshamee));
  XOR stupefiedmclean (.A(kindherschel), .B(dazzlingjerry), .Y(condescendingsatoshi));
  XOR tenderjunior (.A(optimisticvarahamihira), .B(sadjimmy), .Y(jovialhenrietta));
  XOR tenderkilby (.A(compassionatejose), .B(naughtyjangles), .Y(greatmoser));
  XOR thirstyjay (.A(trustingcolden), .B(pensivehailey), .Y(lovingkowalevski));
  XOR thirstyjulieta (.A(confidentbouman), .B(heuristicgagarin), .Y(elatedhedgie));
  XOR thirstypoitras (.A(peacefuljackson), .B(frostyjasmine), .Y(friendlyjenny));
  XOR unruffledjohanna (.A(sleepygypsy), .B(vibranthodgkin), .Y(quizzicalpanini));
  XOR wizardlykerchak (.A(adoringhook), .B(strangekhorana), .Y(kindherschel));
  XOR xenodochiallovelace (.A(cooljackjack), .B(pedantichumbert), .Y(niceclarke));
  XOR youthfulhugo (.A(pedantickhayyam), .B(practicaljubileena), .Y(modestmontalcini));
  XOR youthfulshannon (.A(tenderellis), .B(amazingkermit), .Y(friendlyhamilton));
  XOR youthfulwilbur (.A(confidentbouman), .B(ecstaticsinoussi), .Y(pricelesskalam));
  XOR zealousharry (.A(boldishizaka), .B(joviallehmann), .Y(excitinghoonah));
  XOR zealoushoover (.A(elegantdavinci), .B(competentaustin), .Y(reverentjohn));
  XOR zeniridessa (.A(trustinghades), .B(optimisticvarahamihira), .Y(inspiringisabela));
  assign { y[15], y[7] } = { x[15], x[7] };
  assign agitatedbose = x[6];
  assign blissfulalbattani = x[13];
  assign crankykeldysh = x[10];
  assign eagerpoincare = x[9];
  assign ecstaticsinoussi = x[1];
  assign heuristicchaum = x[12];
  assign infalliblejoy = x[0];
  assign naughtynapier = x[3];
  assign optimisticvarahamihira = x[5];
  assign sleepygypsy = x[11];
  assign sweetimelda = x[8];
  assign unruffledgwen = x[4];
  assign youthfulantonelli = x[14];
  assign youthfulturing = x[2];
  assign y[13] = pricelesskevin;
  assign y[14] = elatedharper;
  assign y[9] = elegantkaa;
  assign y[10] = quirkymendel;
  assign y[11] = dreamygustavo;
  assign y[12] = pedanticmeninsky;
  assign y[8] = sadgould;
  assign y[0] = hopefulhaibt;
  assign y[1] = nicejoshamee;
  assign y[2] = jovialgyro;
  assign y[3] = niceclarke;
  assign y[4] = sharpheffalump;
  assign y[5] = excitinghoonah;
  assign y[6] = elasticborg;
endmodule
